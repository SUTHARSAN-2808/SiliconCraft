module orgate(input x,
          input y,
          output z);
  or org(z,x,y);
endmodule
