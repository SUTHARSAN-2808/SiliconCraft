interface inter;
  
  logic clk;
  logic reset;
  logic d;
  logic [3:0] out;
  
endinterface
