
interface dfff;
  logic reset;
  logic d;
  logic q;
  logic clk;
endinterface
