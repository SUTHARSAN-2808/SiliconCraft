module And(input x,
           input y,
           output z);
  and (z,x,y);
endmodule

