module norgate(input x,
               input y,
               output z);
  nor nor1(z,x,y);
endmodule
