class transaction;
  
  bit clk;
  bit reset;
  bit d;
  reg [3:0]out;
  
endclass
