class transaction;
 rand bit a;
 rand bit b;
 rand bit cin;
  reg sum;
  reg cout;
  
//  constraint 
endclass
