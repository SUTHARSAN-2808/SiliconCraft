class transaction;
  
  rand bit rd;
  bit clk;
  bit reset;
   rand bit [3:0]datain;
  bit [3:0] dataout;
  bit wen;
  bit ren;
  bit full;
  bit empty;
  
endclass
