interface inter;
  logic clk;
  logic reset;
  logic wen;
  logic ren;
  logic [3:0]datain;
  logic [3:0] dataout;
  logic full;
  logic empty;
endinterface
