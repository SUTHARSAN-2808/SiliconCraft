module nand_gate(input x,
                 input y,
                 output z);
  nand (z,x,y);
endmodule
