module Strings;
 string s1="Jai";
  string s2="Akash";
  string s3="Surendhar";
  string s4,s5,s6;
  initial begin
  s4="sutharsan";
  s5="Roja";
    s6="";
    
    $display("s1=%s,s2=%s,s3=%s,s4=%s,s5=%s,s6=%s",s1,s2,s3,s4,s5,s6);
  end
endmodule

