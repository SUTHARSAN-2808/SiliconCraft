interface count_if #(parameter N=2) ;  
logic reset,clk;  
logic [N:0] counter;
endinterface:count_if
